`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.03.2024 12:00:28
// Design Name: 
// Module Name: ACC_MATRIX_MUL_TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module ACC_MATRIX_MUL_TB();
// Inputs
	reg clk;
	reg reset;
	reg [287:0] data_arr;
	reg [287:0] wt_arr;

	// Outputs
	wire [287:0] acc_result1;wire [287:0] acc_result2;wire [287:0] acc_result3;
	wire [287:0] acc_result4;wire [287:0] acc_result5;wire [287:0] acc_result6;
	wire [287:0] acc_result7;wire [287:0] acc_result8;wire [287:0] acc_result9;
	// Instantiate the Unit Under Test (UUT)
	ACC_MATRIX_MULTI dut (
		.clk(clk), 
		.reset(reset), 
		.data_arr(data_arr), 
		.wt_arr(wt_arr), 
		.acc_result1(acc_result1),
		.acc_result2(acc_result2),
		.acc_result3(acc_result3),
		.acc_result4(acc_result4),
		.acc_result5(acc_result5),
		.acc_result6(acc_result6),
		.acc_result7(acc_result7),
		.acc_result8(acc_result8),
		.acc_result9(acc_result9)
	);
always #5 clk = ~clk;
    	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		data_arr <=288'h 000000000000000000000000000000000000000000000000000000000000000000000000;
		wt_arr <=288'h 000000000000000000000000000000000000000000000000000000000000000000000000;
		
		#5
		#10
		reset=0;
		wt_arr<=288'h 404000000000000000000000000000000000000000000000000000000000000000000000;
		data_arr<=288'h 3f8000000000000000000000000000000000000000000000000000000000000000000000;
		
		#10
		wt_arr<=288'h 400000004080000000000000000000000000000000000000000000000000000000000000;
		data_arr<=288'h 3f8000004000000000000000000000000000000000000000000000000000000000000000;
		
		#10
		wt_arr<=288'h 404000003f80000040000000000000000000000000000000000000000000000000000000;
		data_arr<=288'h 3f8000004000000000000000000000000000000000000000000000000000000000000000;

		#10
		wt_arr<=288'h 3f80000040000000408000003f8000000000000000000000000000000000000000000000;
		data_arr<=288'h 3f8000003f8000003f8000003f8000000000000000000000000000000000000000000000;
		
		#10
		wt_arr<=288'h 3f8000003f8000003f8000003f8000003f80000000000000000000000000000000000000;
		data_arr<=288'h 3f8000003f800000404000003f8000003f80000000000000000000000000000000000000;
		
		#10
		wt_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f800000000000000000000000000000;
		data_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f800000000000000000000000000000;
		
		#10
		wt_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000000000000000000000;
		data_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000000000000000000000;
		
		#10
		wt_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000003f80000000000000;
		data_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000003f80000000000000;
		
		#10
		wt_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 3f8000003f8000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 000000003f8000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 000000003f8000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 00000000000000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 00000000000000003f8000003f8000003f8000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 0000000000000000000000003f8000003f8000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 0000000000000000000000003f8000003f8000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 000000000000000000000000000000003f8000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 000000000000000000000000000000003f8000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 00000000000000000000000000000000000000003f8000003f8000003f8000003f800000;
		data_arr<=288'h 00000000000000000000000000000000000000003f8000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 0000000000000000000000000000000000000000000000003f8000003f8000003f800000;
		data_arr<=288'h 0000000000000000000000000000000000000000000000003f8000003f8000003f800000;
		
		#10
		wt_arr<=288'h 000000000000000000000000000000000000000000000000000000003f8000003f800000;
		data_arr<=288'h 000000000000000000000000000000000000000000000000000000003f8000003f800000;
		
		#10
		wt_arr<=288'h 00000000000000000000000000000000000000000000000000000000000000003f800000;
		data_arr<=288'h 00000000000000000000000000000000000000000000000000000000000000003f800000;
		
		#110 $finish;
		
		end
      
endmodule
	
